library ieee;
use ieee.std_logic_1164.all;

entity controlunit_tb is
end controlunit_tb;

architecture TB_ARCHITECTURE of controlunit_tb is
	-- Component declaration of the tested unit
	component controlunit
	port(
		clk_in : in STD_LOGIC;
		reset_in : in STD_LOGIC;
		alu_op_in : in STD_LOGIC_VECTOR(4 downto 0);
		stage_out : out STD_LOGIC_VECTOR(5 downto 0)
	);
	end component;

	-- Stimulus signals
	signal clk_in : STD_LOGIC := '0';
	signal reset_in : STD_LOGIC := '0';
	signal alu_op_in : STD_LOGIC_VECTOR(4 downto 0) := (others => '0');
	signal stage_out : STD_LOGIC_VECTOR(5 downto 0);

	-- Clock period definition
	constant CLK_PERIOD : time := 10 ns;

begin
	-- Unit Under Test port map
	UUT : controlunit
		port map (
			clk_in => clk_in,
			reset_in => reset_in,
			alu_op_in => alu_op_in,
			stage_out => stage_out
		);

	-- Clock signal generation
	clk_process : process
	begin
		clk_in <= '0';
		wait for CLK_PERIOD / 2;
		clk_in <= '1';
		wait for CLK_PERIOD / 2;
	end process;

	-- Stimulus process
	stimulus_process : process
	begin
		-- Initial reset
		reset_in <= '1';
		alu_op_in <= "00000";
		wait for CLK_PERIOD * 2; 

		reset_in <= '0';
		wait for CLK_PERIOD;

		-- Test different ALU operations
		alu_op_in <= "00001";
		wait for CLK_PERIOD * 5;

		alu_op_in <= "00110";
		wait for CLK_PERIOD * 5;

		alu_op_in <= "11111";
		wait for CLK_PERIOD * 5;


		report "Testbench completed successfully";
		wait;
	end process;

end TB_ARCHITECTURE;

configuration TESTBENCH_FOR_controlunit of controlunit_tb is
	for TB_ARCHITECTURE
		for UUT : controlunit
			use entity work.controlunit(behavioral);
		end for;
	end for;
end TESTBENCH_FOR_controlunit;
